--ALU_1BIT Implementation
--By Kenneth Willeford
--This module will take in 2 inputs, a carry in, a control signal, 
-- Given 00 it will send out the 'and' of the inputs.
-- Given 01 it will send out the 'or' of the inputs.
-- Given 10 it will give out the sum of the inputs. 
-- Given 11 it will give out '0'.
-- It will send out the carry out of the sum regardless of signal.
-- All values will be calculated and then a result chosen.
library ieee;
use ieee.std_logic_1164.all;


entity ALU_1BIT is
port(	a,b,cin,sig0,sig1: in std_logic;
		result,cout: out std_logic
);
end ALU_1BIT;

architecture struct of ALU_1BIT is
   component MUX4X1 is
	port(	input1,input2,input3,input4,sig0,sig1: in std_logic;
		result: out std_logic
	);
   end component;
   
   component ORG is
   port( x1,x2: in std_logic;
         y1: out std_logic
	);
   end component;
   component ANDG is
   port( x1,x2: in std_logic;
         y1: out std_logic
	);
   end component;

	component ADD is
	port(	a,b,cin: in std_logic;
			sum,cout: out std_logic
	);
	end component;
	
   signal or_result,and_result,sum_result: std_logic;	
begin

	SUM_RES: ADD  port map (a,b,cin,sum_result,cout);	--	Get Sum and send out Carry Out
	OR_RES:	 ORG  port map (a,b,or_result);				--	Get Or Result
	AND_RES: ANDG port map (a,b,and_result);			--	Get And Result
	Final_Result: MUX4X1 port map (and_result,or_result,sum_result,'0',sig0,sig1,result);	-- Send out result based on signal.
end struct;